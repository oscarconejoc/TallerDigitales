//Oscar Conejo 2020234423

module adder (
    input logic [31:0] A,
    input logic [31:0] B,
    output logic [31:0] out,
);
    
    assign out = A + B;


endmodule